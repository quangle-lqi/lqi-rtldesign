always @(posedge clk)